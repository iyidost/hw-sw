library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity vga_rom_obstacle2 is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(8 downto 0);
      data: out std_logic_vector(15 downto 0)
   );
end vga_rom_obstacle2;

architecture arch of vga_rom_obstacle2 is
   constant ADDR_WIDTH: integer:=9;
   constant DATA_WIDTH: integer:=16;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant obstacle2_ROM: rom_type:=(  -- 2^9-by-16
-- OBSTACLE2 
-- Tile #1
X"0000",X"0000",X"07FF",X"0C00",X"1800",X"3000",X"2000",X"2000",X"3000",X"1800",X"0C00",X"07FF",X"00E0",X"0039",X"000F",X"0030",
-- Tile #2
X"0000",X"0000",X"FFC0",X"0060",X"0030",X"0018",X"0008",X"0008",X"0018",X"0030",X"0060",X"FFC0",X"6000",X"8000",X"E000",X"F800",
-- Tile #3
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"01C0",X"01CF",X"01F8",X"03C0",X"0381",X"07FE",X"0700",X"2F00",
-- Tile #4
X"0000",X"0000",X"0000",X"0001",X"0003",X"0006",X"0006",X"0FE6",X"F026",X"0023",X"0022",X"03E2",X"FC22",X"0022",X"0021",X"00C0",
-- Tile #5
X"0000",X"0000",X"FFFF",X"8000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"C000",
-- Tile #6
X"0000",X"0000",X"F800",X"0C00",X"0600",X"0300",X"0100",X"0100",X"0300",X"FFFC",X"0004",X"0004",X"0004",X"000C",X"0018",X"0020",
-- Sprite empty 110 
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0FFF",X"0FFF",X"0C20",X"0C20",X"0C20",
-- Sprite empty 111
X"0000",X"0000",X"0000",X"0000",X"07FF",X"1C00",X"1800",X"1800",X"1800",X"1800",X"1800",X"D800",X"D800",X"5800",X"5FFF",X"4FFF",


-- Tile #7
X"0030",X"000C",X"0003",X"0000",X"0000",X"0180",X"0180",X"0383",X"031E",X"03FC",X"0780",X"0E00",X"0C00",X"0C00",X"0C00",X"0C00",
-- Tile #8
X"0780",X"01F0",X"803E",X"E00F",X"3001",X"6000",X"CC00",X"1300",X"10C0",X"1060",X"1020",X"1020",X"1020",X"1020",X"1020",X"1020",
-- Tile #9
X"3F00",X"3AFF",X"5200",X"D200",X"527F",X"1780",X"1400",X"247F",X"4C80",X"8FFF",X"B000",X"A000",X"A000",X"A000",X"A000",X"A000",
-- Tile #10
X"7F00",X"8400",X"0400",X"0C00",X"F400",X"0400",X"7C00",X"8401",X"0406",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
-- Tile #11
X"4000",X"4000",X"4000",X"4000",X"4000",X"4000",X"C000",X"8000",X"0000",X"FEFF",X"0300",X"0080",X"0060",X"0020",X"0020",X"0020",
-- Tile #12
X"0040",X"0080",X"0100",X"0100",X"0108",X"0208",X"0218",X"0218",X"0218",X"E3A8",X"20E8",X"2008",X"1008",X"1008",X"1008",X"1008",
-- Sprite empty 110 
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0FFF",X"0FFF",X"0C20",X"0C20",X"0C20",
-- Sprite empty 111
X"0000",X"0000",X"0000",X"0000",X"07FF",X"1C00",X"1800",X"1800",X"1800",X"1800",X"1800",X"D800",X"D800",X"5800",X"5FFF",X"4FFF",


-- Tile #13
X"0C00",X"0C00",X"0C00",X"0E00",X"0780",X"03FC",X"031E",X"0383",X"0180",X"0180",X"0000",X"0000",X"0003",X"000C",X"0030",X"0030",
-- Tile #14
X"1020",X"1020",X"1020",X"1020",X"1020",X"1060",X"10C0",X"1300",X"CC00",X"6000",X"3001",X"E00F",X"803E",X"01F0",X"0780",X"F800",
-- Tile #15
X"A000",X"A000",X"A000",X"A000",X"B000",X"8FFF",X"4C80",X"247F",X"1400",X"1780",X"527F",X"D200",X"5200",X"3AFF",X"3F00",X"2F00",
-- Tile #16
X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0406",X"8401",X"7C00",X"0400",X"F400",X"0C00",X"0400",X"8400",X"7F00",X"00C0",
-- Tile #17
X"0020",X"0020",X"0060",X"0080",X"0300",X"FEFF",X"0000",X"8000",X"C000",X"4000",X"4000",X"4000",X"4000",X"4000",X"4000",X"C000",
-- Tile #18
X"1008",X"1008",X"1008",X"2008",X"20E8",X"E3A8",X"0218",X"0218",X"0218",X"0208",X"0108",X"0100",X"0100",X"0080",X"0040",X"0020",
-- Sprite empty 110 
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0FFF",X"0FFF",X"0C20",X"0C20",X"0C20",
-- Sprite empty 111
X"0000",X"0000",X"0000",X"0000",X"07FF",X"1C00",X"1800",X"1800",X"1800",X"1800",X"1800",X"D800",X"D800",X"5800",X"5FFF",X"4FFF",



-- Tile #19
X"000F",X"0039",X"00E0",X"07FF",X"0C00",X"1800",X"3000",X"2000",X"2000",X"3000",X"1800",X"0C00",X"07FF",X"0000",X"0000",X"0000",
-- Tile #20
X"E000",X"8000",X"6000",X"FFC0",X"0060",X"0030",X"0018",X"0008",X"0008",X"0018",X"0030",X"0060",X"FFC0",X"0000",X"0000",X"0000",
-- Tile #21
X"0700",X"07FE",X"0381",X"03C0",X"01F8",X"01CF",X"01C0",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
-- Tile #22
X"0021",X"0022",X"FC22",X"03E2",X"0022",X"0023",X"F026",X"0FE6",X"0006",X"0006",X"0003",X"0001",X"0000",X"0000",X"0000",X"0000",
-- Tile #23
X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"8000",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #24
X"0018",X"000C",X"0004",X"0004",X"0004",X"FFFC",X"0300",X"0100",X"0100",X"0300",X"0600",X"0C00",X"F800",X"0000",X"0000",X"0000",







others => X"0000");
signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= obstacle2_ROM(to_integer(unsigned(addr_reg)));
end arch;




