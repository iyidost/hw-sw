library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity vga_rom_obstacle3_inv is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(8 downto 0);
      data: out std_logic_vector(15 downto 0)
   );
end vga_rom_obstacle3_inv;

architecture arch of vga_rom_obstacle3_inv is
   constant ADDR_WIDTH: integer:=9;
   constant DATA_WIDTH: integer:=16;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant obstacle3_inv_ROM: rom_type:=(  -- 2^9-by-16
-- OBSTACLE3 
-- Tile #1
X"0000",X"0000",X"003F",X"003F",X"0FE0",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0921",X"0926",
-- Tile #2
X"0000",X"0000",X"FFFF",X"FFFF",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"FFFF",X"0000",
-- Tile #3
X"0000",X"3FFF",X"C000",X"FFFF",X"0800",X"0800",X"0800",X"0871",X"0800",X"0800",X"0807",X"081C",X"0862",X"0B81",X"FE01",X"31C0",
-- Tile #4
X"0000",X"FFFF",X"0000",X"FFFF",X"0000",X"4000",X"4000",X"C000",X"4000",X"4000",X"FFC0",X"00B8",X"0086",X"0081",X"8080",X"C100",
-- Tile #5
X"0000",X"FFFF",X"0000",X"FFFF",X"0800",X"0E00",X"0980",X"0880",X"0D43",X"0D4C",X"0AA0",X"0AA0",X"09E0",X"8860",X"FFFF",X"4060",
-- Tile #6
X"0000",X"FFFF",X"0000",X"FFFF",X"0380",X"0E00",X"3000",X"C000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"1000",
-- Tile #7
X"0000",X"FFC0",X"0070",X"FFFF",X"6808",X"7808",X"787F",X"784D",X"784D",X"784D",X"784D",X"787F",X"580C",X"380C",X"FFFF",X"3400",
-- Tile #8
X"0000",X"0000",X"0000",X"F000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"F000",X"1000",


-- Tile #9
X"0938",X"07E0",X"0040",X"0040",X"0041",X"0043",X"0042",X"0044",X"004C",X"0040",X"0043",X"00C6",X"0048",X"0070",X"0040",X"0040",
-- Tile #10
X"4018",X"4063",X"819F",X"8670",X"1D80",X"6600",X"8400",X"0400",X"4400",X"C400",X"0400",X"0400",X"0C00",X"0C00",X"0400",X"0400",
-- Tile #11
X"C030",X"000E",X"E001",X"1FC0",X"0000",X"0000",X"0000",X"001F",X"0010",X"0020",X"0030",X"0018",X"000C",X"0007",X"0000",X"0000",
-- Tile #12
X"6100",X"310F",X"DAF0",X"2C00",X"05F0",X"000F",X"0000",X"8000",X"8000",X"FFFE",X"0422",X"FFFE",X"8000",X"0000",X"0000",X"0000",
-- Tile #13
X"A118",X"1107",X"1900",X"0900",X"0700",X"E180",X"1FE0",X"0018",X"3FFF",X"2000",X"2000",X"1000",X"1000",X"1000",X"1000",X"1000",
-- Tile #14
X"1003",X"007C",X"E7C0",X"1800",X"1600",X"1300",X"10C1",X"1033",X"F00A",X"0804",X"0804",X"0804",X"0804",X"07FF",X"0000",X"0000",
-- Tile #15
X"CC00",X"1400",X"247F",X"6F80",X"4800",X"8807",X"0438",X"00E0",X"0700",X"0400",X"0400",X"0400",X"FFFF",X"0100",X"0100",X"0100",
-- Tile #16
X"1000",X"1000",X"D000",X"3C00",X"1C00",X"E000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"FFFF",X"8101",X"8101",X"8101",


-- Tile #17
X"0040",X"0070",X"0048",X"00C6",X"0043",X"0040",X"004C",X"0044",X"0042",X"0043",X"0041",X"0040",X"0040",X"07E0",X"0938",X"0926",
-- Tile #18
X"0400",X"0C00",X"0C00",X"0444",X"0482",X"C4BA",X"44BA",X"0482",X"84FE",X"6600",X"1D80",X"8670",X"819F",X"4063",X"4018",X"0000",
-- Tile #19
X"006C",X"0182",X"0201",X"0100",X"0100",X"0100",X"0100",X"0181",X"00C2",X"0024",X"0018",X"1FC0",X"E001",X"000E",X"C030",X"31C0",
-- Tile #20
X"0000",X"0000",X"8000",X"8000",X"8000",X"8000",X"8000",X"8000",X"0000",X"0007",X"03F0",X"2E00",X"DAF0",X"310F",X"6100",X"C100",
-- Tile #21
X"1000",X"1000",X"1000",X"1000",X"2000",X"2000",X"3FFF",X"0018",X"1FE0",X"E180",X"0700",X"0900",X"1900",X"1107",X"A118",X"4060",
-- Tile #22
X"0000",X"07FF",X"0804",X"0804",X"0804",X"0804",X"F00A",X"1033",X"10C1",X"1300",X"1600",X"1800",X"E7C0",X"007C",X"1003",X"1000",
-- Tile #23
X"0100",X"0100",X"FFFF",X"0400",X"0400",X"0400",X"0700",X"00E0",X"0438",X"8807",X"4800",X"6F80",X"247F",X"1400",X"CC00",X"3400",
-- Tile #24
X"8101",X"8101",X"FFFF",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"E000",X"1C00",X"3C00",X"D000",X"1000",X"1000",X"1000",


-- Tile #25
X"0921",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0920",X"0FE0",X"003F",X"003F",X"0000",X"0000",X"0000",
-- Tile #26
X"FFFF",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"103F",X"1000",X"1000",X"1000",X"FFFF",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #27
X"FE01",X"0B81",X"0862",X"081C",X"0807",X"0800",X"0800",X"C871",X"0800",X"0800",X"0800",X"FFFF",X"C000",X"3FFF",X"0000",X"0000",
-- Tile #28
X"8080",X"0081",X"0086",X"00B8",X"FFC0",X"4000",X"4000",X"C000",X"4000",X"4000",X"0000",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #29
X"FFFF",X"8860",X"09E0",X"0AA0",X"0AA0",X"0D4C",X"0D43",X"0880",X"0980",X"0E00",X"0800",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #30
X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"C000",X"3000",X"0E00",X"0380",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #31
X"FFFF",X"380C",X"580C",X"787F",X"784D",X"784D",X"784D",X"784D",X"787F",X"7808",X"6808",X"FFFF",X"0070",X"FFC0",X"0000",X"0000",
-- Tile #32
X"F000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"1000",X"F000",X"0000",X"0000",X"0000",X"0000",


others => X"0000");
signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= obstacle3_inv_ROM(to_integer(unsigned(addr_reg)));
end arch;




