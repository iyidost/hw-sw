library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity vga_rom_obstacle3_inv is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(8 downto 0);
      data: out std_logic_vector(15 downto 0)
   );
end vga_rom_obstacle3_inv;

architecture arch of vga_rom_obstacle3_inv is
   constant ADDR_WIDTH: integer:=9;
   constant DATA_WIDTH: integer:=16;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant obstacle3_inv_ROM: rom_type:=(  -- 2^9-by-16
-- OBSTACLE3 
-- Tile #1
X"0000",X"0000",X"0000",X"0000",X"001F",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DE",X"06D9",
-- Tile #2
X"0000",X"0000",X"0000",X"0000",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"0000",X"FFFF",
-- Tile #3
X"0000",X"0000",X"3FFF",X"0000",X"F7FF",X"F7FF",X"F7FF",X"F78E",X"F7FF",X"F7FF",X"F7F8",X"F7E3",X"F79D",X"F47E",X"01FE",X"CE3F",
-- Tile #4
X"0000",X"0000",X"FFFF",X"0000",X"FFFF",X"BFFF",X"BFFF",X"3FFF",X"BFFF",X"BFFF",X"003F",X"FF47",X"FF79",X"FF7E",X"7F7F",X"3EFF",
-- Tile #5
X"0000",X"0000",X"FFFF",X"0000",X"F7FF",X"F1FF",X"F67F",X"F77F",X"F2BC",X"F2B3",X"F55F",X"F55F",X"F61F",X"779F",X"0000",X"BF9F",
-- Tile #6
X"0000",X"0000",X"FFFF",X"0000",X"FC7F",X"F1FF",X"CFFF",X"3FFF",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"0000",X"EFFF",
-- Tile #7
X"0000",X"0000",X"FF80",X"0000",X"97F7",X"87F7",X"8780",X"87B2",X"87B2",X"87B2",X"87B2",X"8780",X"A7F3",X"C7F3",X"0000",X"CBFF",
-- Tile #8
X"0000",X"0000",X"0000",X"0000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"0000",X"E000",


-- Tile #9
X"06C7",X"001F",X"003F",X"003F",X"003E",X"003C",X"003D",X"003B",X"0033",X"003F",X"003C",X"0039",X"0037",X"000F",X"003F",X"003F",
-- Tile #10
X"BFE7",X"BF9C",X"7E60",X"798F",X"E27F",X"99FF",X"7BFF",X"FBFF",X"BBFF",X"3BFF",X"FBFF",X"FBFF",X"F3FF",X"F3FF",X"FBFF",X"FBFF",
-- Tile #11
X"3FCF",X"FFF1",X"1FFE",X"E03F",X"FFFF",X"FFFF",X"FFFF",X"FFE0",X"FFEF",X"FFDF",X"FFCF",X"FFE7",X"FFF3",X"FFF8",X"FFFF",X"FFFF",
-- Tile #12
X"9EFF",X"CEF0",X"250F",X"D3FF",X"FA0F",X"FFF0",X"FFFF",X"7FFF",X"7FFF",X"0001",X"FBDD",X"0001",X"7FFF",X"FFFF",X"FFFF",X"FFFF",
-- Tile #13
X"5EE7",X"EEF8",X"E6FF",X"F6FF",X"F8FF",X"1E7F",X"E01F",X"FFE7",X"C000",X"DFFF",X"DFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",
-- Tile #14
X"EFFC",X"FF83",X"183F",X"E7FF",X"E9FF",X"ECFF",X"EF3E",X"EFCC",X"0FF5",X"F7FB",X"F7FB",X"F7FB",X"F7FB",X"F800",X"FFFF",X"FFFF",
-- Tile #15
X"33FF",X"EBFF",X"DB80",X"907F",X"B7FF",X"77F8",X"FBC7",X"FF1F",X"F8FF",X"FBFF",X"FBFF",X"FBFF",X"0000",X"FEFF",X"FEFF",X"FEFF",
-- Tile #16
X"E000",X"E000",X"2000",X"C000",X"E000",X"0000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"0000",X"7EFE",X"7EFE",X"7EFE",


-- Tile #17
X"003F",X"000F",X"0037",X"0039",X"003C",X"003F",X"0033",X"003B",X"003D",X"003C",X"003E",X"003F",X"003F",X"001F",X"06C7",X"06D9",
-- Tile #18
X"FBFF",X"F3FF",X"F3FF",X"FBBB",X"FB7D",X"3B45",X"BB45",X"FB7D",X"7B01",X"99FF",X"E27F",X"798F",X"7E60",X"BF9C",X"BFE7",X"FFFF",
-- Tile #19
X"FF93",X"FE7D",X"FDFE",X"FEFF",X"FEFF",X"FEFF",X"FEFF",X"FE7E",X"FF3D",X"FFDB",X"FFE7",X"E03F",X"1FFE",X"FFF1",X"3FCF",X"CE3F",
-- Tile #20
X"FFFF",X"FFFF",X"7FFF",X"7FFF",X"7FFF",X"7FFF",X"7FFF",X"7FFF",X"FFFF",X"FFF8",X"FC0F",X"D1FF",X"250F",X"CEF0",X"9EFF",X"3EFF",
-- Tile #21
X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"DFFF",X"DFFF",X"C000",X"FFE7",X"E01F",X"1E7F",X"F8FF",X"F6FF",X"E6FF",X"EEF8",X"5EE7",X"BF9F",
-- Tile #22
X"FFFF",X"F800",X"F7FB",X"F7FB",X"F7FB",X"F7FB",X"0FF5",X"EFCC",X"EF3E",X"ECFF",X"E9FF",X"E7FF",X"183F",X"FF83",X"EFFC",X"EFFF",
-- Tile #23
X"FEFF",X"FEFF",X"0000",X"FBFF",X"FBFF",X"FBFF",X"F8FF",X"FF1F",X"FBC7",X"77F8",X"B7FF",X"907F",X"DB80",X"EBFF",X"33FF",X"CBFF",
-- Tile #24
X"7EFE",X"7EFE",X"0000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"0000",X"E000",X"C000",X"2000",X"E000",X"E000",X"E000",


-- Tile #25
X"06DE",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"06DF",X"001F",X"0000",X"0000",X"0000",X"0000",X"0000",
-- Tile #26
X"0000",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFFF",X"EFC0",X"EFFF",X"EFFF",X"EFFF",X"0000",X"0000",X"0000",X"0000",X"0000",
-- Tile #27
X"01FE",X"F47E",X"F79D",X"F7E3",X"F7F8",X"F7FF",X"F7FF",X"378E",X"F7FF",X"F7FF",X"F7FF",X"0000",X"3FFF",X"0000",X"0000",X"0000",
-- Tile #28
X"7F7F",X"FF7E",X"FF79",X"FF47",X"003F",X"BFFF",X"BFFF",X"3FFF",X"BFFF",X"BFFF",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #29
X"0000",X"779F",X"F61F",X"F55F",X"F55F",X"F2B3",X"F2BC",X"F77F",X"F67F",X"F1FF",X"F7FF",X"0000",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #30
X"0000",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"FFFF",X"3FFF",X"CFFF",X"F1FF",X"FC7F",X"0000",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #31
X"0000",X"C7F3",X"A7F3",X"8780",X"87B2",X"87B2",X"87B2",X"87B2",X"8780",X"87F7",X"97F7",X"0000",X"FF80",X"0000",X"0000",X"0000",
-- Tile #32
X"0000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"E000",X"0000",X"0000",X"0000",X"0000",X"0000",


others => X"0000");
signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= obstacle3_inv_ROM(to_integer(unsigned(addr_reg)));
end arch;




