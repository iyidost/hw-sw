library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity vga_rom_obstacle3_layer1 is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(8 downto 0);
      data: out std_logic_vector(15 downto 0)
   );
end vga_rom_obstacle3_layer1;

architecture arch of vga_rom_obstacle3_layer1 is
   constant ADDR_WIDTH: integer:=9;
   constant DATA_WIDTH: integer:=16;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant obstacle3_ROM: rom_type:=(  -- 2^9-by-16
-- OBSTACLE 3 layer 1
-- Tile #1
X"0000",X"0000",X"0000",X"000F",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"000F",X"0008",
-- Tile #2
X"0000",X"03FF",X"0E00",X"FFFF",X"1016",X"101E",X"FE1E",X"B21E",X"B21E",X"B21E",X"B21E",X"FE1E",X"301A",X"301C",X"FFFF",X"002C",
-- Tile #3
X"0000",X"FFFF",X"0000",X"FFFF",X"01C0",X"0070",X"000C",X"0003",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0008",
-- Tile #4
X"0000",X"FFFF",X"0000",X"FFFF",X"0010",X"0070",X"0190",X"0110",X"C2B0",X"32B0",X"0550",X"0550",X"0790",X"0611",X"FFFF",X"0602",
-- Tile #5
X"0000",X"FFFF",X"0000",X"FFFF",X"0000",X"0002",X"0002",X"0003",X"0002",X"0002",X"03FF",X"1D00",X"6100",X"8100",X"0101",X"0083",
-- Tile #6
X"0000",X"FFFC",X"0003",X"FFFF",X"0010",X"0010",X"0010",X"8E10",X"0010",X"0010",X"E010",X"3810",X"4610",X"81D0",X"807F",X"038C",
-- Tile #7
X"0000",X"0000",X"FFFF",X"FFFF",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"FFFF",X"0000",
-- Tile #8
X"0000",X"0000",X"FC00",X"FC00",X"07F0",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"8490",X"6490",



-- Tile #9
X"0008",X"0008",X"000B",X"003C",X"0038",X"0007",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"FFFF",X"8081",X"8081",X"8081",
-- Tile #10
X"0033",X"0028",X"FE24",X"01F6",X"0012",X"E011",X"1C20",X"0700",X"00E0",X"0020",X"0020",X"0020",X"FFFF",X"0080",X"0080",X"0080",
-- Tile #11
X"C008",X"3E00",X"03E7",X"0018",X"0068",X"00C8",X"8308",X"CC08",X"500F",X"2010",X"2010",X"2010",X"2010",X"FFE0",X"0000",X"0000",
-- Tile #12
X"1885",X"E088",X"0098",X"0090",X"00E0",X"0187",X"07F8",X"1800",X"FFFC",X"0004",X"0004",X"0008",X"0008",X"0008",X"0008",X"0008",
-- Tile #13
X"0086",X"F08C",X"0F5B",X"0034",X"0FA0",X"F000",X"0000",X"0001",X"0001",X"7FFF",X"4420",X"7FFF",X"0001",X"0000",X"0000",X"0000",
-- Tile #14
X"0C03",X"7000",X"8007",X"03F8",X"0000",X"0000",X"0000",X"F800",X"0800",X"0400",X"0C00",X"1800",X"3000",X"E000",X"0000",X"0000",
-- Tile #15
X"1802",X"C602",X"F981",X"0E61",X"01B8",X"0066",X"0021",X"0020",X"0022",X"0023",X"0020",X"0020",X"0030",X"0030",X"0020",X"0020",
-- Tile #16
X"1C90",X"07E0",X"0200",X"0200",X"8200",X"C200",X"4200",X"2200",X"3200",X"0200",X"C200",X"6300",X"1200",X"0E00",X"0200",X"0200",


-- Tile #17
X"8081",X"8081",X"FFFF",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0007",X"0038",X"003C",X"000B",X"0008",X"0008",X"0008",
-- Tile #18
X"0080",X"0080",X"FFFF",X"0020",X"0020",X"0020",X"00E0",X"0700",X"1C20",X"E011",X"0012",X"01F6",X"FE24",X"0028",X"0033",X"002C",
-- Tile #19
X"0000",X"FFE0",X"2010",X"2010",X"2010",X"2010",X"500F",X"CC08",X"8308",X"00C8",X"0068",X"0018",X"03E7",X"3E00",X"C008",X"0008",
-- Tile #20
X"0008",X"0008",X"0008",X"0008",X"0004",X"0004",X"FFFC",X"1800",X"07F8",X"0187",X"00E0",X"0090",X"0098",X"E088",X"1885",X"0602",
-- Tile #21
X"0000",X"0000",X"0001",X"0001",X"0001",X"0001",X"0001",X"0001",X"0000",X"E000",X"0FC0",X"0074",X"0F5B",X"F08C",X"0086",X"0083",
-- Tile #22
X"3600",X"4180",X"8040",X"0080",X"0080",X"0080",X"0080",X"8180",X"4300",X"2400",X"1800",X"03F8",X"8007",X"7000",X"0C03",X"038C",
-- Tile #23
X"0020",X"0030",X"0030",X"2220",X"4120",X"5D23",X"5D22",X"4120",X"7F21",X"0066",X"01B8",X"0E61",X"F981",X"C602",X"1802",X"0000",
-- Tile #24
X"0200",X"0E00",X"1200",X"6300",X"C200",X"0200",X"3200",X"2200",X"4200",X"C200",X"8200",X"0200",X"0200",X"07E0",X"1C90",X"6490",

-- Tile #25
X"000F",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"000F",X"0000",X"0000",X"0000",X"0000",
-- Tile #26
X"FFFF",X"301C",X"301A",X"FE1E",X"B21E",X"B21E",X"B21E",X"B21E",X"FE1E",X"101E",X"1016",X"FFFF",X"0E00",X"03FF",X"0000",X"0000",
-- Tile #27
X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0003",X"000C",X"0070",X"01C0",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #28
X"FFFF",X"0611",X"0790",X"0550",X"0550",X"32B0",X"C2B0",X"0110",X"0190",X"0070",X"0010",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #29
X"0101",X"8100",X"6100",X"1D00",X"03FF",X"0002",X"0002",X"0003",X"0002",X"0002",X"0000",X"FFFF",X"0000",X"FFFF",X"0000",X"0000",
-- Tile #30
X"807F",X"81D0",X"4610",X"3810",X"E010",X"0010",X"0010",X"8E13",X"0010",X"0010",X"0010",X"FFFF",X"0003",X"FFFC",X"0000",X"0000",
-- Tile #31
X"FFFF",X"0008",X"0008",X"0008",X"0008",X"0008",X"0008",X"FC08",X"0008",X"0008",X"0008",X"FFFF",X"FFFF",X"0000",X"0000",X"0000",
-- Tile #32
X"8490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"0490",X"07F0",X"FC00",X"FC00",X"0000",X"0000",X"0000",

others => X"0000");
signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= obstacle3_ROM(to_integer(unsigned(addr_reg)));
end arch;




