library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity vga_rom_sprites is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(8 downto 0);
      data: out std_logic_vector(15 downto 0)
   );
end vga_rom_sprites;

architecture arch of vga_rom_sprites is
   constant ADDR_WIDTH: integer:=9;
   constant DATA_WIDTH: integer:=16;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant HEX2LED_ROM: rom_type:=(  -- 2^9-by-16
----------------------------------------------------------
-- Memory data for the car pics (current one tile only) --
----------------------------------------------------------
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0FFF",X"8000",
X"0000",X"07FF",X"C000",X"0000",X"3800",X"E000",X"0000",X"1C00",
X"7000",X"0000",X"3000",X"6000",X"0000",X"1800",X"3000",X"0000",
X"3000",X"6000",X"0000",X"1800",X"3000",X"0000",X"3000",X"6000",
X"0000",X"1800",X"3000",X"0000",X"3000",X"6000",X"0000",X"1800",
X"3000",X"0000",X"3000",X"6000",X"0000",X"1800",X"3000",X"0000",
X"3000",X"6000",X"0FFF",X"D800",X"3000",X"0000",X"3000",X"6000",
X"0FFF",X"D800",X"3000",X"0000",X"3000",X"6000",X"0C20",X"5800",
X"3000",X"0000",X"3FFF",X"E000",X"0C20",X"5FFF",X"F00F",X"FFFF",
X"9FFF",X"C000",X"0C20",X"4FFF",X"E018",X"0000",X"4068",X"0000",
X"0C20",X"4078",X"0030",X"0000",X"2068",X"0000",X"0C20",X"C078",
X"0060",X"0000",X"1068",X"0000",X"0C21",X"806C",X"00C0",X"0000",
X"0868",X"0000",X"0C22",X"006E",X"0180",X"0000",X"0468",X"0000",
X"0C24",X"0066",X"0300",X"0000",X"0668",X"0000",X"0C28",X"0067",
X"0600",X"0000",X"02C8",X"0000",X"0C28",X"0063",X"0C00",X"0000",
X"018B",X"FFF8",X"0C28",X"0063",X"9800",X"0000",X"008A",X"1218",
X"0C30",X"0061",X"F000",X"07FE",X"004B",X"FFF8",X"0C30",X"007F",
X"FFFF",X"F803",X"802A",X"1218",X"0C38",X"3FC0",X"0000",X"0000",
X"E03E",X"1218",X"0C27",X"E000",X"0001",X"FFE0",X"3802",X"1218",
X"0C27",X"0000",X"0006",X"0037",X"0E02",X"1218",X"0C38",X"0000",
X"0008",X"C013",X"E382",X"1218",X"0C20",X"0000",X"0008",X"C011",
X"38E2",X"1218",X"0C20",X"0000",X"000F",X"C011",X"0C3A",X"1218",
X"0C20",X"0000",X"0008",X"C011",X"38E2",X"1218",X"0C38",X"0000",
X"0008",X"C013",X"E382",X"1218",X"0C27",X"0000",X"0006",X"0037",
X"0E02",X"1218",X"0C27",X"E000",X"0001",X"FFE0",X"3802",X"1218",
X"0C38",X"3FC0",X"0000",X"0000",X"E03E",X"1218",X"0C30",X"007F",
X"FFFF",X"F803",X"802A",X"1218",X"0C30",X"0061",X"F000",X"07FE",
X"004A",X"1218",X"0C28",X"0063",X"9800",X"0000",X"008A",X"1218",
X"0C28",X"0063",X"0C00",X"0000",X"018B",X"FFF8",X"0C28",X"0067",
X"0600",X"0000",X"02CA",X"1218",X"0C24",X"0066",X"0300",X"0000",
X"066B",X"FFF8",X"0C22",X"006E",X"0180",X"0000",X"0468",X"0000",
X"0C21",X"806C",X"00C0",X"0000",X"0868",X"0000",X"0C20",X"C078",
X"0060",X"0000",X"1068",X"0000",X"0C20",X"4078",X"0030",X"0000",
X"2068",X"0000",X"0C20",X"4FFF",X"E018",X"0000",X"4068",X"0000",
X"0C20",X"5FFF",X"F00F",X"FFFF",X"9FFF",X"C000",X"0C20",X"5800",
X"3000",X"0000",X"3FFF",X"E000",X"0FFF",X"D800",X"3000",X"0000",
X"3000",X"6000",X"0FFF",X"D800",X"3000",X"0000",X"3000",X"6000",
X"0000",X"1800",X"3000",X"0000",X"3000",X"6000",X"0000",X"1800",
X"3000",X"0000",X"3000",X"6000",X"0000",X"1800",X"3000",X"0000",
X"3000",X"6000",X"0000",X"1800",X"3000",X"0000",X"3000",X"6000",
X"0000",X"1800",X"3000",X"0000",X"3000",X"6000",X"0000",X"1C00",
X"7000",X"0000",X"3000",X"6000",X"0000",X"07FF",X"C000",X"0000",
X"3800",X"E000",X"0000",X"0000",X"0000",X"0000",X"0FFF",X"8000",
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
others => X"0000");
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= HEX2LED_ROM(to_integer(unsigned(addr_reg)));
end arch;